* series resonant bandpass filter
V1 0 1 ac 1 dc 0
Rs 1 2 100
R1 2 3 375
C2 2 0 20e-12
C1 3 4 33.0e-15
L1 4 0 30e-3
*Rl 4 0 50
*Cf 1 5 0.1e-12
*Cq 5 0 8.4e-12
*Rf 1 5 10
*Rl 1 0 1e5

.control
ac lin 100000 4.900e6 5.163e6
write test.raw all
